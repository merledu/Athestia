`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/29/2025 03:13:55 PM
// Design Name: 
// Module Name: verifyTop_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module verifyTop_tb(


module verifyTop_tb;
    // Define parameters inside the testbench
    parameter int PK_SIZE = 20736;  // 2592 bytes
    parameter int MSG_MAX_SIZE = 25624; // Maximum message size
    parameter int SIG_SIZE = 37016;  // 4627 bytes
    parameter int CTX_SIZE = 2032;
    
    
    logic clk;
    logic rst;
    logic [PK_SIZE-1:0] pk;  
    logic [MSG_MAX_SIZE-1:0] M;
    logic [SIG_SIZE-1:0] sigma;  
    logic valid;  // Assume 'valid' is an output from the DUT
    logic initial_start;
    logic [CTX_SIZE-1:0]ctx;

    // Instantiate the Device Under Test (DUT)
    VerifyTop #(
        .PK_SIZE(PK_SIZE),  //  2592  bytes
        .MSG_MAX_SIZE(MSG_MAX_SIZE),    // Maximum message size (adjustable)
        .SIG_SIZE(SIG_SIZE)  
    ) dut (
        .clk(clk),
        .rst(rst),
        .pk(pk),
        .M(M),
        .sigma(sigma),
        .valid(valid),
        .start(initial_start),
        .ctx(ctx)
    );

    // Clock generation (Toggle every 0.5 time units)

    // Testbench sequence
    initial begin
        clk = 1; // Initialize clock 
        rst = 1'b1;
        pk = 0;
        M = 0;
        sigma = 0;
        ctx = 0;
        initial_start = 1'b0;

        #1;  // Wait for some time before finishing the simulation
        rst=1'b0;
        initial_start = 1'b1;
             
//               big endian reverse
                   ctx = 2032'hEF4F61C539431EBF5BA1C912F40AAC18C2719EB8E9F26E07DA503947E684FAE7AD21DECC243682F5EFCFF7761B613D3B3E7915FE462326FDE059EAE809D6D8D7A7E265D22CE0F48BEEA8C919FAF7EC7812FE096D6EFBA08AFBE0EBCA4C9AEC18F620CF38FC6B0F5E858A0F9D5A0C02E86D72D50BCD6B69AB41DBD74BF4293F54BCB022DA28B37BA7EFABE7E4EB022FEFDD025DD9C4E14B8BB624F62193C36A5B4ABBE1A9E927C0B9F62E1B218384BF3FABE86DF1CC658FDB65972304BD5A132C418B9A30218605B642A3E395C529073264B775AB55788FE42B05435204BCFC9B1AEFE0F7EA8F1D25E2B7AE2882FA163C8FF19F05E568D6C8FCB5041B42B3;
                   pk = 20736'hE6BEC0F78BE5941B0C42A54CEB8A3AB62CF0A59495C90837647202E361E7480F123A0B4B3F4698657EE88A14CB13CE45FE28791F09FCC4E24584FC11778E6513BA6B659166923B020A8E99E8F3D2D3A2D5C2619B192500D5B6BF22E580C892E3DC2D02AB9FEE2448D9E2B2EE2783E563301731AFCD98DC913C6F697D1D99D32582FFF20BC91354CA32D2436A82D5CB7B96834150D9E3AA4A79EF3A55634AD6745035ACBBAD68983A9A766B73EFA346C2734D0D5D6D88497974D85A3719867996D303F417AB26C1A359EB60952D3930344B829A8C767E9D1ED2361D0157CA27E3BBC8C1BBD5C7112E9E7525A44D6875A03C914EE2CF5622F2D66BFE08DA799CF99587FF0D4E0A4509C4CE22322F22FDA680A14DFF362E02CB4F1E73CB1800A9D447F39883C5598B0721ECF1DEAD9D7AA09D077C89AB520CDDA5C9CF9A2EA7B3A68BF3355FB4709EAA533773C353BC5D07AB4E1AE820976F2D9A9FCC84CD7032514D107346D68C2C45E0D2EEE1ADC3FB011E3FD079E3830414DE1FC412786EB65FEF537AC7FAD48A3B7E2A054184CFBAA17C007098AF1C9D1B866A8533B24C1FD480679C06C2CFEA049991BF41C8FBAFFB093D1F16EFFB2FBE2701056A58A500A72DEDCD34AFEC303B902691D33D13273D68F4A5DD419EB2F86FF495EC2A9E4CADD951DBF56F2E6D1F9BE3487366DA21697BD9DDC18EF62512904E6D49CDC4FF601BE26BE69968F60A005A8AFE87E60919D8A5383BAFED66A5151D17B634EB2EBD36B6FE9265C2B96022845CDD9A5594C834670C0104C8D563489F0129B289AC88BAC746F0A3F8AF37E8D95259BF1E1CE77FBA690FAB5ADCDD2B64FA709C3EA40BCB801FAB828ADFD96B46A51096712A0A5C5F87084B9FFC42C9C8F02326D17CA2DCE50160CE4BC58B7789242DB8A3B1A0A627B0D39811CE99487AEBB6E65C00F794FA2DC5921C16F244FEB2EA952C4847B4E44B21433833ACAF0E20CEB7793932DBB2DB7274C522BE0D5935E822109422A4E6B15F15CC2BE3D001B523A6D8B6419AC71619B6C844E5FAC92A53C25F88095727AA130016951B9E96326B9B598ABD09D9024D2957D37861F67DD2D8843D0DEF74F9C9752D5C5D9A7705E5C505A887FAA6B360211BE88F0C2C0344A8DE7B27E0D8C85B590682DE22F1C173C387C101A7393461AA1F7DD21C43A61AD5524D67A01E2E13D2F565FBAEB892CCBA4E3798AC9B38CAA40584E055C4B4C5CEF11C6323516FE27F7C851A2C7ACEE5539A773C9EF32EFFC617B304EB4E71B134EF71F00F7462D20ADB090B1DE55EF366033645BB65D79DC49E45DD6C27B4C0CC4D1DE84F4D01D2DC755975690263DB4201F6642CCD3C71AF8065623EA92F780729A969C959897DA6F2B3E2508BE6827D6F864A70A7F8F6F3B3A058BC638089313840C24AC5AC96A1196AD510EBBECC0BCB5ADC19E59DD51FEA3984AF3FEB33B742D62D2EC01950037C59B67F99F59A29886428978713B183D792CB9AF8EA03ABAF29CD8038115B8DC68E59DE2A6780C7DD7454395C009175AE43D79B5F4A5EED130C065E9280520246D6AAB12180DEE721FCB5D6AE90D65B80BE8A30D339589E9C82DB010BECE1DA8AA18118C010D4086D357053748F40180DDA0877ACCF68692865D87EBF0D69416A5F7AD77DA39568B9A32D1C1FFE99309231CFA7674AE23113B91FE36D8225D294202156CD9DA95D6D0D06B73B50990DF82CCE407B1ECA14DF861AEF399D923E4F5C5E3EE2CD2661C050CBDF1511F3A6B3E8FD1B5662380450DCD6D673A11998A46824338BD9D68E50215ABA2757834DE3A570654CDCBD57F67AB777761D5D2694E7D808A747409D7598514BB93A46C9F1ABD3247C0A6AA16424B3EBAFC1C8FD43AC5C5CE2EFB5CC85D52463C696E406F8F2A2E0F4A3DD2794BA1CDEC4850856A30D1FCAB77F0DD689F29775D3E295FAD65B4074E30B069AC0418D384CA7A1DE498E9097AC993D2FCE34400DA4C9FC392F7EC12F619058764C6CC283B45C63A6DAD5C1B549168504FE834F99CA2A129AF7922064A761FE6128ADBCA32DC0F4F96283B0A45573DCB6067FFED2782D3C304F9B25083AA551B0588664728E8A1FEC4F920EF7EA8554B27F0695F904B80A1A3054B37A745B3CE0D6BECA3554042C0142E189FC9A7FE127766755F216D6D736322A7A7AE3BEEB19497F9DF304B9EAB1F310FD343E4ED0A751BD78A87EFF34D20A5D4C78F5B096C63C436D29D147426892B9188921E4A450493390848BC7C7255EF1937EB17903FCDE48C6CF331D7148C37AE07C8D9DDB55F2063D63F46B98ABE2E4A13C752B2639A82382F37E58A239CF9E65863A412AF40A806EDDCC78436E96C377993C3181277CF8C1A2BF25B4F5551BD9E9094A0C79850DE4C9692600EA2F0CFB404713ABF827D58972400892F37CB6000E83E4FA89420F592836739D2A49A9B87E4678D700C0225E4C297FA1EF1C3E5745383C858C6A9CC980D33D38F220D1085D45DE8E8E893E43AAAECE58A3E6F8960E054A0651BA70B592686734401CD45253E85697A2431D2BC246B3D1EE432DE7410ED6633FEFF4C44658F3D9281E341ED4BB6950E0CD6BB47D1A296344D650D451E0A9E3437E2F59C6A77F7C9C2B84D90D6DF81612952381795F75329EACAF79F3F2F81FE8916EC6638DDFF11313A185DD8D3FBBB64AFC85B7CC52F6129F106247A875C7D00479EF51B1ABAD38FE909F9AF9F8D86FBA2C740A3454B7854D8AA16720DEB55D2CC414733357B0EB9A5A7F321552C5B788FF23387F430693EAB3A8087B8F7552DBBFECCB31B315FC33A6AF28197F35F20609062B135B7229CF96D0345436B769662B3A38BF6461EF6BF7FB879DB3860838630F804A69EE5A14B34B1FB4612C1F06908A46C034823CFC26549240ACF731DA480526C866E6BE2004B94A4DFD9D778771BF8732DC871C2C9A832A6873447D31F67191B924AA77FB040E8E0EBF8EC5FF6D58F4FD02EFF656A8CF95C229C513A1FC90743EFF8A6E3CF0F235F2002A22AC3F1D127689CD5F7804C2E417F9DFD1D87BD89DFA5C9CAB21517A09030965E76AE84893A0FDFB644086B7B162ADD5DC15D51FCCE553CDAF738C8D72E9D53BFA334567358533CC58297BC2E4BD65182AD1D27FA802823EBEFD2034E3D5560494C4D34D30F6621C02DE005A582A1990B497A7D70B1D770AB0C7860968C2AE80A2B6E9EC1D9524CF386B2B1FFAB6DD2A4DEE883BF4814337043CACC66B69750C24B710DB161B65566395897D211BBE05986D29ABA05A58457B2C56B7CD110AA79EC1A3842C9FCA7F6AC3831B5F8BB9A4FD11C26D82E7BD59AF12698487C6EF3FBB4361C09BD090508C6EE7349C0553C7F217DF1BA20ABB0A477996BA5A09DC27E3DB0120A9106A68C044F7080DFC23F336598ECA5A3C25DD298B034D45965E2BB7A67E1D7CDB4373E5511406C23CAC51B9444B5F6E90602E3E02EB6B015420E0A8B0A1EAF8C599E06F75C3B1DEB01DD80D376037B769653D96F7F14512D6337B624AC70DC45CE19D1BFF5F5B8EFE6DF01AB6A5C0CC32B70500EBBAAE9F23BFD5F77D5E8FC79311BEF8053390FA6F4A74C26B510797D7252C7E07650EC0BAFE1B91E31917825D7ABF198033A0F02517147CD20977721F106614B964C8D13FEAF76C68F0EA;
                  M = 25624'hFFCB5B1267B32866626139C37A5CC724B1C7B67ABB44F50D7384B1774BEF8D44175BED314BBE63EF382A968EB888B640C4FE90955B8AFFBBD54D9EE302B11A73D4F5AC1F6E96D8F263C64190AD6754EBCD70B24C5FF7E98C5C325CFE1F80EC870F23B9C3DC97D12D269D3194496E0D6DF9B31592FECD14DC0B1FC23B3ADAD3E3D9B9808AAD900E369E8526C1C55443ED25EE056B6A5A89410FDDB7BCD496F34BCA4EBA8FED82BF68A5DFF378A75216B7DCD5164BD467787E2F3E7BD0D852610891DAF77799B3FFA22E9DC68A67109ABCC600E0FF80A77662D53C60AF07EF8F527DEAE7CC5A9F1D28D5731C37A1EE171EA4BE09D8716288E96395A15D53509A3F0D730C7C29CD6227E2B8290C8A3FC1E724410A49E5B6E11B62FD69C5FDBFD485D8DD292DE19AF5D65BE2F5B9397B5F24D3BA381245515A5692F11A2C649C2A22E3A333AD1594068A4C33ED03C127E2E69E44F14287C23F8782D39AEF7FC872BFB7D2D59547B10F3FB4AEC5116357956A0F348E1FAAE79B2164AC2B42F9160A83C12E4BEE514C9EED35B28ED8FC2D232A3D30E04B3A5214D037B4309B85CC469DA34250350CA718C295A0EAF858C32436880005C835BF486F1A7AB69C1C0367686BF135BADDEE1E95171EB599671B777490F91285C77D67E3F9E11B91F07BA69139818D678D6A599AE16FB11709AF07FE02420C22F0E2A0ED8951C0FCD38DA49B772460E68E10E626A078A358CC4FDA4AD91C8EAD6F84A057E19FDD3CA95DC754CA15A0E54E2170F25CE681783E482039777622B6FFF72CF3830905EE32A97C42B14F8DB7AFF4FBB8AB9C5188022818987EA4C5323A1055D3E9AD62451C82BFB2693EC7EFBA698A827A6A0A63A5A3F05BF06C6F8EE44A07A0FABACD0292B69C29DC9E1FC36029DE151942B8D006F22D45BC0754B01331CD1F3627F4009B88F0C3CDE18606832CFAC78D5974A291369A088C88458B62EC16ABD1008C3934DE799152F403246B27C18F0C8C22B9BC2B8DFF8CEC7413426461E1CADB35839FC193AFE0E34F9D33759C65C6B57ED6C95DEEA5728CAD4769654FED93225A8FF13EF04BF872D8D9DBF0CC16500F4D8CE58A176DEC8F1113144C457A94620A111B0C7387C533DD578415CA82C096F65A18C207080AECA3612CDD37AC2D5E4579E6BAFB439BC5C7B2ADC0E9D6C58F527D55EA62D15A01062F69125BE8FC302926D0519C059AB3BF52FA555B4A03CC9C9D8AB95742FB731EE4B3CCDA896ADFB67C96C20674F34CE3A22B10D704A5BC2B9C75BD5D42D9E72A5D32B752CED836E81B9FDEB440C628AA3DD6B517EB9B1A3EF7A03D13AC8173A3AF98A8413BFA14C9F528BB65C607EBD64D13206C24D03FC218785A2E9A223B9A2B3B05A81EE66E43C1EB22C3DFB478EFB467C59860077FDE58E629C39FE62ED2EC213A8B0243B867A4DCAB38AD7CE263006B79335DA23924BC264F37BCABA3DABC4FD6BE7AECEC71AE5EF4845C4630DB03C6C3346DFB7549E715CFDCF380AAF939D07C5EA623E8137E0884FEAEB5C875F57433F6E86F6DC1DA8CD6641D107D2EB3FA4B8BCAD235DFDDAFB56576769B324D59E67F4CB411C963BB83194D83F66D8B564BB36A3CAB223E531838B9084A64F1A317C329FDE1FEE981280F4E1B9259B948D91F2AE7C811AEC441F99CD8105B701F28A96C32438D754DCAE8139BD422C1BE7F712E2A3909DB051565BCE8611071CD9E2EF3E8ED86044BA9DC1DDFFD12F01E37DE589E2C45E61FCE661DDED18DECB97746FDA52FD8D1F96CE2805CECFB0802759DB083B8D2A05848D31A866926791CF06367B7154AEE5E0D5F324AC48933D25E1B6834DD6801A5A5A45C5CBE4A8F4668646B889350EC2AAE517658A05693BEA048284EBD453F8862C21171EE92A0C2CFEBE2601DAA3E0D2E3D858BF2A8054F109DBB762241892225E326D13F7B3C1CB0B388B47433A1F5091A1F7FC0B395B9BDC26050D72AA08E62BF3B39846DCEB30169DA3F2050DBDCFCC56C07220962714E6C137C1AEC448612FA52B4F867719C4B6C7E56D855996DE7845311BD996B595CC9EB175952981424542D25FD26E49553D0BBB58A0B99F8D3A595969833C8798EF9582F7C5943F9D4693284287470C19FBDBDEDDDB6CE502FF244B3BC027CF18BB49603CDB519FA8DC1E120D915D05F35D4F6DB75DB9BD82A07FF89158F3DD1ED40F874DD6CF3EAA4C3601CD5AE761A22E57DE80BA07CB018BED9C6B58FE4FD840F32981C5B81C9E00C36B17A7F037C90E5672F1154C64CC4485B1E932D3414DF6297C57BDEFDC664B407FE6ACB3599BB5D35D028B5EB3049E5D4D4FF6236B3D722D217E83D00B2E7A1CB5C4CC7E2F913C26335F763EB2977677C960A29C6017E542647F91DB17D5D82E887E98FE38102DAC03CFE00BB7436A8A080C069A8BEDACADEF8A09B00F611E5D8757A6440E783FB932F6889027E98B210507C30BCF3DA2AAC1FB0EBE067DACA2B192746F9D268B8FDC5D5795650C75F60ED8BAF79E128E49A50B72037981A2C549D5EE95651B93EE8C332F61D60D45C57518BF2DC2B5149F042ACA81A478165ABA925B8F2DE090E344DC6B6AE32C6397B5BC8E50D2750284C14F913A51023A041CC4B743B1B6979477CBE8F659A9ABE7B722DBF7F9B588458FC6CDDE5F56923292574E1E652FE5FF24E9E9068C1C3B1793B9733E36321A574C61B3FAF8B9452129B653F25B8D72973CDCD30FDC71B9739BA64AA5D363FC503CF6D1F36BFAF66BA4B7ECD5C838BC0636EBF1696F0A7ACAB8405F527E9F4DB5B9F3B564BB7F2B41D6675B2494D3BB62EA346EF77292F1327C074B2B9BA3FD056A272BC473575AC7B0AF8307BF5635D484FC683A305643170282E8A423FFB6227A45BA6DA7E6FF92E99736C31FE97325C166A69F4BB2D513D414C1E06EA693C0E9508D69ABD82CAE0CC550991F7007191FC2D2CD5916E6B770968993250F24330375E9BF5C1979F939F89276623C04641DA8D0ABD3D667C279D5E9054E9988FD911D95A99647BCF648D98350846045449225757C3E886F2D0E1735863074BAA07FA4D554966ACDC5FBDA52FA43074E1990A47329140CBF18AE689B7F1236C5D42EE2E0DF8AF0AE2757BF80643574E9F6C92BF59BF1818C62E5CCA63DCF4EB3B5147ECB50266E8E9FF65BC1648C5AD3398E94B5F64139E2AD667DF9CE4A705808FBCB4FB6B999C06A9D5595A5C027E69AE97CAF3A98CD73EA9C2DF9B874B05585F3B868C10B2C8FE4C45B58FB944CED4E976ED4DDC12D703E47651A9BA017E5DCF01FA207BF158FCCFCBA664D7488465F30AB2115EB87B4D6482A799601E444BC657BFB849AE58F71DF17D106B722C9CF2ECB5AF4E6DFF1785ADBBF94ABE9BB0875A9E7F89CC1C45B2BBF36C3A6AE1F2560BA7746995FC5857A8329BF25FAC5F55CD8911D4AC1325CF6FFC937A92DC1BCCC8A23F162746F15E4527E19A8052530E94176CE1CF1DA9F882A4F99869DEC5CB17CF29BC6D482E8697B38F84328B4F1CA984E67B7039FCABF94794824D59F566621583B02896A14BE9E6491C8E24C5F755DDEEE4F8495BDDD37EC225B4AB393EBD28221C079EF312E39A9189EFDF1CD4819D2D706A116E18BAA5DDAAD37B973DAC0B5F6502A9EFB6E9DC005DB7D1EDF361EEA4177EC9D4ACBA096161C0493F670354DCE480B7D2D7AD76868E101160E9B8EA48E5D780BEE336B2ABF9488DF69F9D985A63F40873AA1BCC690842469CA8A877A9D60159908295F9ADCE0BD98E207FE7F078B7FDF5AF779DCA0A17B5A1F0150251D1E4209E4307D7CDFA5BA49F423D49885B5524F1AA82F95E638E866BE058BCB80887BD3C5F48AD70E030FA54D2FE87CCCE2C469BF111A64EEAC13BB5816BEDA29EEC96BA7F0C2912A8B3117A87A58C6406B99DB31221C6F7E16F519E0DF8EE744258B5E668CD4CC10333F33DFF2CC74434D6AEC7CD3A907D259ED910BB8A05B0C59C372FEFA6FC396DDCAFDE2D88F8B4A70D69364927A708C738C0C9F33B06792E437862F497548EDA745AF08AB14F9CA62469AD20CE669DF52F67B6E5324531D636B0EA1095C00FB8DB5BD5CCB67D16E92423CED258585FDDDA6DC5309DA9A82E281A5401658C106459F5457390D03FB151CDC10E775F7DDE500C3528FADF1A31B2A6A49B28148397126A796312EB4C092E13DFD0E79AB7C99C76B05856E8697ADA13C0E92CA3883C4929FB0CE61ACB64C02BFAE7FF4A4918EFDBFFB2642B402A00FE88FF2A63DD8A8AA286BE9EAAE381AB4B982BEE827A90C9A8FA51A4D6D81EE9D10CE792CC395D4E6F5D5CC38B7944F77D071893153B7E84F83582688BE6B3CA68D5CD9EFCEFDE113BDC7E251DCC3D2FB55926CFBF8BD3958E629A96B7F4C289A9925BB6ABA6FB8D28065739BD59672BF752B332BFE40ADC01370F995547594619F57C8B7087830E5E98A6B9339AD835FB6E9F654190C9C4877EB473966138E0AC101FC7DDDCBA70CEA4D3263D51A9675FDA9EE6A8F405892BB703F1D21077FC60C60C227B10;
//                  27672'hFFCB5B1267B32866626139C37A5CC724B1C7B67ABB44F50D7384B1774BEF8D44175BED314BBE63EF382A968EB888B640C4FE90955B8AFFBBD54D9EE302B11A73D4F5AC1F6E96D8F263C64190AD6754EBCD70B24C5FF7E98C5C325CFE1F80EC870F23B9C3DC97D12D269D3194496E0D6DF9B31592FECD14DC0B1FC23B3ADAD3E3D9B9808AAD900E369E8526C1C55443ED25EE056B6A5A89410FDDB7BCD496F34BCA4EBA8FED82BF68A5DFF378A75216B7DCD5164BD467787E2F3E7BD0D852610891DAF77799B3FFA22E9DC68A67109ABCC600E0FF80A77662D53C60AF07EF8F527DEAE7CC5A9F1D28D5731C37A1EE171EA4BE09D8716288E96395A15D53509A3F0D730C7C29CD6227E2B8290C8A3FC1E724410A49E5B6E11B62FD69C5FDBFD485D8DD292DE19AF5D65BE2F5B9397B5F24D3BA381245515A5692F11A2C649C2A22E3A333AD1594068A4C33ED03C127E2E69E44F14287C23F8782D39AEF7FC872BFB7D2D59547B10F3FB4AEC5116357956A0F348E1FAAE79B2164AC2B42F9160A83C12E4BEE514C9EED35B28ED8FC2D232A3D30E04B3A5214D037B4309B85CC469DA34250350CA718C295A0EAF858C32436880005C835BF486F1A7AB69C1C0367686BF135BADDEE1E95171EB599671B777490F91285C77D67E3F9E11B91F07BA69139818D678D6A599AE16FB11709AF07FE02420C22F0E2A0ED8951C0FCD38DA49B772460E68E10E626A078A358CC4FDA4AD91C8EAD6F84A057E19FDD3CA95DC754CA15A0E54E2170F25CE681783E482039777622B6FFF72CF3830905EE32A97C42B14F8DB7AFF4FBB8AB9C5188022818987EA4C5323A1055D3E9AD62451C82BFB2693EC7EFBA698A827A6A0A63A5A3F05BF06C6F8EE44A07A0FABACD0292B69C29DC9E1FC36029DE151942B8D006F22D45BC0754B01331CD1F3627F4009B88F0C3CDE18606832CFAC78D5974A291369A088C88458B62EC16ABD1008C3934DE799152F403246B27C18F0C8C22B9BC2B8DFF8CEC7413426461E1CADB35839FC193AFE0E34F9D33759C65C6B57ED6C95DEEA5728CAD4769654FED93225A8FF13EF04BF872D8D9DBF0CC16500F4D8CE58A176DEC8F1113144C457A94620A111B0C7387C533DD578415CA82C096F65A18C207080AECA3612CDD37AC2D5E4579E6BAFB439BC5C7B2ADC0E9D6C58F527D55EA62D15A01062F69125BE8FC302926D0519C059AB3BF52FA555B4A03CC9C9D8AB95742FB731EE4B3CCDA896ADFB67C96C20674F34CE3A22B10D704A5BC2B9C75BD5D42D9E72A5D32B752CED836E81B9FDEB440C628AA3DD6B517EB9B1A3EF7A03D13AC8173A3AF98A8413BFA14C9F528BB65C607EBD64D13206C24D03FC218785A2E9A223B9A2B3B05A81EE66E43C1EB22C3DFB478EFB467C59860077FDE58E629C39FE62ED2EC213A8B0243B867A4DCAB38AD7CE263006B79335DA23924BC264F37BCABA3DABC4FD6BE7AECEC71AE5EF4845C4630DB03C6C3346DFB7549E715CFDCF380AAF939D07C5EA623E8137E0884FEAEB5C875F57433F6E86F6DC1DA8CD6641D107D2EB3FA4B8BCAD235DFDDAFB56576769B324D59E67F4CB411C963BB83194D83F66D8B564BB36A3CAB223E531838B9084A64F1A317C329FDE1FEE981280F4E1B9259B948D91F2AE7C811AEC441F99CD8105B701F28A96C32438D754DCAE8139BD422C1BE7F712E2A3909DB051565BCE8611071CD9E2EF3E8ED86044BA9DC1DDFFD12F01E37DE589E2C45E61FCE661DDED18DECB97746FDA52FD8D1F96CE2805CECFB0802759DB083B8D2A05848D31A866926791CF06367B7154AEE5E0D5F324AC48933D25E1B6834DD6801A5A5A45C5CBE4A8F4668646B889350EC2AAE517658A05693BEA048284EBD453F8862C21171EE92A0C2CFEBE2601DAA3E0D2E3D858BF2A8054F109DBB762241892225E326D13F7B3C1CB0B388B47433A1F5091A1F7FC0B395B9BDC26050D72AA08E62BF3B39846DCEB30169DA3F2050DBDCFCC56C07220962714E6C137C1AEC448612FA52B4F867719C4B6C7E56D855996DE7845311BD996B595CC9EB175952981424542D25FD26E49553D0BBB58A0B99F8D3A595969833C8798EF9582F7C5943F9D4693284287470C19FBDBDEDDDB6CE502FF244B3BC027CF18BB49603CDB519FA8DC1E120D915D05F35D4F6DB75DB9BD82A07FF89158F3DD1ED40F874DD6CF3EAA4C3601CD5AE761A22E57DE80BA07CB018BED9C6B58FE4FD840F32981C5B81C9E00C36B17A7F037C90E5672F1154C64CC4485B1E932D3414DF6297C57BDEFDC664B407FE6ACB3599BB5D35D028B5EB3049E5D4D4FF6236B3D722D217E83D00B2E7A1CB5C4CC7E2F913C26335F763EB2977677C960A29C6017E542647F91DB17D5D82E887E98FE38102DAC03CFE00BB7436A8A080C069A8BEDACADEF8A09B00F611E5D8757A6440E783FB932F6889027E98B210507C30BCF3DA2AAC1FB0EBE067DACA2B192746F9D268B8FDC5D5795650C75F60ED8BAF79E128E49A50B72037981A2C549D5EE95651B93EE8C332F61D60D45C57518BF2DC2B5149F042ACA81A478165ABA925B8F2DE090E344DC6B6AE32C6397B5BC8E50D2750284C14F913A51023A041CC4B743B1B6979477CBE8F659A9ABE7B722DBF7F9B588458FC6CDDE5F56923292574E1E652FE5FF24E9E9068C1C3B1793B9733E36321A574C61B3FAF8B9452129B653F25B8D72973CDCD30FDC71B9739BA64AA5D363FC503CF6D1F36BFAF66BA4B7ECD5C838BC0636EBF1696F0A7ACAB8405F527E9F4DB5B9F3B564BB7F2B41D6675B2494D3BB62EA346EF77292F1327C074B2B9BA3FD056A272BC473575AC7B0AF8307BF5635D484FC683A305643170282E8A423FFB6227A45BA6DA7E6FF92E99736C31FE97325C166A69F4BB2D513D414C1E06EA693C0E9508D69ABD82CAE0CC550991F7007191FC2D2CD5916E6B770968993250F24330375E9BF5C1979F939F89276623C04641DA8D0ABD3D667C279D5E9054E9988FD911D95A99647BCF648D98350846045449225757C3E886F2D0E1735863074BAA07FA4D554966ACDC5FBDA52FA43074E1990A47329140CBF18AE689B7F1236C5D42EE2E0DF8AF0AE2757BF80643574E9F6C92BF59BF1818C62E5CCA63DCF4EB3B5147ECB50266E8E9FF65BC1648C5AD3398E94B5F64139E2AD667DF9CE4A705808FBCB4FB6B999C06A9D5595A5C027E69AE97CAF3A98CD73EA9C2DF9B874B05585F3B868C10B2C8FE4C45B58FB944CED4E976ED4DDC12D703E47651A9BA017E5DCF01FA207BF158FCCFCBA664D7488465F30AB2115EB87B4D6482A799601E444BC657BFB849AE58F71DF17D106B722C9CF2ECB5AF4E6DFF1785ADBBF94ABE9BB0875A9E7F89CC1C45B2BBF36C3A6AE1F2560BA7746995FC5857A8329BF25FAC5F55CD8911D4AC1325CF6FFC937A92DC1BCCC8A23F162746F15E4527E19A8052530E94176CE1CF1DA9F882A4F99869DEC5CB17CF29BC6D482E8697B38F84328B4F1CA984E67B7039FCABF94794824D59F566621583B02896A14BE9E6491C8E24C5F755DDEEE4F8495BDDD37EC225B4AB393EBD28221C079EF312E39A9189EFDF1CD4819D2D706A116E18BAA5DDAAD37B973DAC0B5F6502A9EFB6E9DC005DB7D1EDF361EEA4177EC9D4ACBA096161C0493F670354DCE480B7D2D7AD76868E101160E9B8EA48E5D780BEE336B2ABF9488DF69F9D985A63F40873AA1BCC690842469CA8A877A9D60159908295F9ADCE0BD98E207FE7F078B7FDF5AF779DCA0A17B5A1F0150251D1E4209E4307D7CDFA5BA49F423D49885B5524F1AA82F95E638E866BE058BCB80887BD3C5F48AD70E030FA54D2FE87CCCE2C469BF111A64EEAC13BB5816BEDA29EEC96BA7F0C2912A8B3117A87A58C6406B99DB31221C6F7E16F519E0DF8EE744258B5E668CD4CC10333F33DFF2CC74434D6AEC7CD3A907D259ED910BB8A05B0C59C372FEFA6FC396DDCAFDE2D88F8B4A70D69364927A708C738C0C9F33B06792E437862F497548EDA745AF08AB14F9CA62469AD20CE669DF52F67B6E5324531D636B0EA1095C00FB8DB5BD5CCB67D16E92423CED258585FDDDA6DC5309DA9A82E281A5401658C106459F5457390D03FB151CDC10E775F7DDE500C3528FADF1A31B2A6A49B28148397126A796312EB4C092E13DFD0E79AB7C99C76B05856E8697ADA13C0E92CA3883C4929FB0CE61ACB64C02BFAE7FF4A4918EFDBFFB2642B402A00FE88FF2A63DD8A8AA286BE9EAAE381AB4B982BEE827A90C9A8FA51A4D6D81EE9D10CE792CC395D4E6F5D5CC38B7944F77D071893153B7E84F83582688BE6B3CA68D5CD9EFCEFDE113BDC7E251DCC3D2FB55926CFBF8BD3958E629A96B7F4C289A9925BB6ABA6FB8D28065739BD59672BF752B332BFE40ADC01370F995547594619F57C8B7087830E5E98A6B9339AD835FB6E9F654190C9C4877EB473966138E0AC101FC7DDDCBA70CEA4D3263D51A9675FDA9EE6A8F405892BB703F1D21077FC60C60C227B10EF4F61C539431EBF5BA1C912F40AAC18C2719EB8E9F26E07DA503947E684FAE7AD21DECC243682F5EFCFF7761B613D3B3E7915FE462326FDE059EAE809D6D8D7A7E265D22CE0F48BEEA8C919FAF7EC7812FE096D6EFBA08AFBE0EBCA4C9AEC18F620CF38FC6B0F5E858A0F9D5A0C02E86D72D50BCD6B69AB41DBD74BF4293F54BCB022DA28B37BA7EFABE7E4EB022FEFDD025DD9C4E14B8BB624F62193C36A5B4ABBE1A9E927C0B9F62E1B218384BF3FABE86DF1CC658FDB65972304BD5A132C418B9A30218605B642A3E395C529073264B775AB55788FE42B05435204BCFC9B1AEFE0F7EA8F1D25E2B7AE2882FA163C8FF19F05E568D6C8FCB5041B42B3FE00;
               
//               athstia python direct input
                sigma = 37016'hc883516adee991a12ab7e5fc58fc426438baaa45fcc13b5e222380b85a5c0b0fb8dc8aac10e4cfc921bc7cd18e18a379a539e8cf3fe48f352c43f6aa22c320989f16a7d41b582bdf35531a18cd0345a312dcf86b076e7213247afcbddd4942381b97d981502e4de5668e1e3ef86fa65b3e20e88212aa657b9507dc519fcbd5411a952d8a54518434d10c8d811c7ca871c5fe2932e495c0567abeac9221b9a42924601f0aa9abc1071a1e86321839c7b89abeb0df520d35c22aadfeb35c166dced57b7ed857aff1f49aa1286840ada3ef34663e4559b290ae408ad0c8284084daa1b27444eecc54948af4f738c68f92ed7ea99118ad8b8b9e9976cba8daef9236b28c6151e0ff931166aebf417104427d0e3ec52f33a61ae2cdeab50a182172a50f94581d567b709e9c1e47fcce492885d99c4aee94355bdd8ae2a665f5c86141cffc3ad947083c6388a822e059aa4100f99ef2b73dfbd30ae9f58205b473b77de96d4f68a3a2b4d03f45f22eb4f50481cf80cd2b7ae60d3edac42644a95b4e1782ef4701855b3bab0ba3ff1a2993ec86dba723bfb699d56f1d6678a4189b9d197d2c715737ac557e3c91c94ffad0b37cd2911680d6637a6ddb7e6a3aa62f4fe3a49502753d511b7ddf9c9322be6fd7e9c8fef40c89b50ee3b72fcab674062f5f44072fd867af9fe3d733c17c519c64291c5ddab18306dd5aecebb3b4db3948fc1d3c9429fbcf39cf0e4bbb7ca7602fe64b9bff29c075e3bc5d952b41fee0b8fd73e0fde3d10e5d9cd21dacf15a68c04f7d10bc1c79257e99f89caf8803fbe6fa8f6569e2cf2dcb52c502794d4f4434fd905304d67f00532dacdc148c8e28c0003926a05f234358ff3ebf6a5d467a898661bacd00d06dd2181eec190e6600d60c4f597f3244d2da6c0bed495203c1cd2cb29e8e1e9999444a800fccbf9dde2c902ee9b3fe22abc0cbf464130f43bb4eb01cdb94b8c91f59ab7da8c0b44e8034d6b49776d4b7364fb209ad6a29fc7ada13a38eb5f43e2f917352286004c909c19dbe7d2707aacf4ecf623a85154608a6d345e3086ac53abaca86c46aec94d751cae8020b2f73b9ed9961afd4682407b107fee23fd2ee0a72fea20a0c01ed6f91dc36f8ce216c8f14738b72f7189cf0bf05030e1e428efbcdda957ba0e7f3a1c770e0d3f0f49487984fd024892ddc1b77de81e52477a8af8065c6817cb2eac763fb498799936569cb9a75b8d6cf7392a4863c7e8fc4345c2ff52aa0d0004bb7370fd188d5a2d79a7f82f8cae209361afcc2d094c5b70af3d355fa1eb75287d87bbee38f618c12e50a74b7948243c5a016f17a956dc960c77ad99e7c48a6432f4ffe5263d8f4394b8252486dbd47aa92fa2f902a063d3bbce2569d5cec09812882e87f60b1c0ad4da54f7ce62756f27db3dc4e4c78fe1e7e947a94aa3c04b0836c576d536572723a5ea12ccc5de9329dcb988268796e66327666aeaf6f21084d42060b4528a43da96a77c35b46c568efdfd4fd715719b5cd025b7335a67e9978f0af5dda895672bd77213fc60aa6d23141c20077a2044e26b465c03e476409778093f38203d6ef7d066e6a9f4d7c7ce0ea3e0120cc173318dac3ab9c844df1faca3abedc5ec5f87c4ec4faf2867f11477982d7ec4ef2bfdee4e7891e4c5fb873ceed9d161be0c2b8243c4e3a82975e80b8cfed52e1ebbcf896768d331e8a9533ed655637907a5af009faa6be2cb0862b6c98c148b25cc8a9612001c500043e579774a8b4b6ceed219ae9b729bd502e9b15c4b95faea817dbee92d99fad7e231acd60ad4d5793a429e1ca43578d35de0da661c659e7954beb5e97d522fd41dc6846625d3bf006dacfe503d3bb549ad641149f1b7cf98961c93adc2580e241dbcef17d9e7b61ee5a19dc106bd11fc84ff565f49f853a861a8c5837d95c26888aeda1b5adf66d15b1e1297939374b96265363ed9901fb034f87f1a42d8eda6f2924fa8ee3de50398086009907663863f93c509bcfb1ba68c53107ff503ebae2ead2b00577c283a79c32f5461b744bc6c512dbe058d512627425a6b0c3d68f0dcbf8beacea39a51a6eff464a32106ea05875a6f5370ed6dfb1ceae6ca3288509fb24870ed4086a34d4257a05d75bd2f7d94775af2a2c05f0de79605289d03b9b92719b118c060c2e9abe6a26cec59040662ca0f45e9be16096d9adfd6983815ac4636732af0648545b57b267f54931cb9b8d0571819ecbfc338618a560ef39240ff4c33d79eec160cbdcc1061a042b85ac0d053cb013383b868ce63f2e9690c8526f8e438de07d58fbc8e3aac636df4462a43eaacd31686027f711ebbd7187987661d6fad9531e4abba24176ae3833d00ffa0c14e50e61dd5b83edb91a597964182e9700821c5495657bdb88f7765eb7bd209f5b633ba8b658c3f3de3d63e94c4eefe84054d85978f4c01b6f13a86d73a677a211d87356c83a55afc3733af5739f3719b7f7d9aa2c677aa0068eb7ce4a58a6e9eb71df5b1123b04b4436ed18797818973af0e32ab8f34041899de1b4e87ce86b32042cfc89b3bed71f24982ef7855a9efa1ca6eca9463081c0a039203c57621ec6dd322318fd14a1cad324a705faf90f411013b4669cb388f7fd43cc59b5eefb2e16f57f8ad5b464e152968b984fcec86325bad6f8e996bdbdd8c03bf11ed7aa9704b82c9500666a3e10bce19bcde499580fdccdb979af707734c1adfb9db4785c9acc0f65f9aeb1b090ef2029566c2eca3e0743e206d781dc939772cbb75ccc5967b56e62702d4ccc73605fd2c6e9da18ce9c108315f3b2d7e5b8b2ada85e63569325cb7205cc0c5b0117a3e3d7770971c1cfbfa9e2da4acc82916da2819f5aefc99a2bf2f564c4885864d9f3329b9d029b7abc0385a0f21637bd5f75e04dbc8f1f5d92eaf4b723c4932c222a0512a8c33f06313091f8ffd186695e006059f792120fc1669f32083bec262a93517af1083eee14752482f7f3dd52739680a0282e13c6203d8c4220c8f53e7ce6624c122349005e4657854b6cff4f8e6ea2cd3156e290021cdaeb760be2ff34c4f4e8ff46c9138c5b55242e9fd355fc5556c4dd211514772fe90bfb6521a9ec0764ee6664cf103e8cb3ae2119565a938bd0e3503eb98d904cf422dd4f6b957f865b5851f9a130c982fdc51a1eb5d6992bc195e84d3d009974cd4ff042db8106e8b3d07de94f7323b454cf4422e92f0c621f5c8146a0cf9692e279ef78c1142a8a2b3589a6d0833ec31be1edf16bc810b15df671f61d116dc70587ce1549d8631f2559d0406a1189903ca73c263dc4d87facecdbdee1d62a8cfc5b9a2600e7305d44733fe25c56ad4a175f1ef16ba689640eada4d0b396d426a0eb4e40850f5f8b15eebc450f4cd0010c69c460eccead862225537b6ee4e053d5c245d8b38f6610b4e1877e2a70f406a203d52cf6c9e227da1a4d817d78f079d9b04c4e80b10d5b870ae4b908fc9c38850d29d3e1413659defd75e55b1fea868ef7c49ffc43e855974083050042b4d72d915c924ae83e671f92c2bdb2ed23dc9b34832c9eded134a107ed321a42f46ed99007834907a1ea4e9c37a18528dc9bd23db7371af48ce1d9184ce4a8a82309507122de7667e0bd40a11c66d86124a4d48e182331c613e18def7b5372348295763e3412247a9d8b142d9ed707426211a49e70d48af13975773066565ce3472716ed2413431f0a1bc36deb5a784c306a29ee1bee261f51f2e97f1f06efc57b985f56ca0365f47a196c48eaefb83ebc1027fe2132bd2db7dc0f9e557a5f535ddb48eca41bc9e01656d3e4513d5968b072d64c30eea5e72065d33d5c6465e5b8aa53068ff9566902a9f1373b366ed1e5a9cdc3499f540825d7bb5a5cb2e40ecd09bd693ef9f021ebe346a71d166220a36971936b6fb04cfe37f4b2e2fdab3094d03c9a0f5d8ad1433369426fd352278903dcdc31ba41b7e981236bf53a830a67060d7586cc5d0a5bf622b297122c746884c101c051c97592204108f470459b22c328d77eec93bb0601d8d8608002874517efbbc9ef6127c48e0b39778731aa2dbefdff93c9bfd47a13aa189c31d2c1ffd64a267c2ceb4dbadaaed1656e97e4cbfa374e762ab18676cf5f7c24f8e67b470bbf83a08a1c2047ecc478dbd8c1d3f19a2f10d79c0895383148b6bd1346d359591389df84084d166f24a005333cfb1a26ecea248ab18e4233f9d3d83b49253cfaf666e2db49e65e66b43b8c41942a6c4dff4100c64d9da5ae48b2284d87e4cb9997e640e7d653d0a658bf14486376c9db6c2ac27b0e560a92b958a20ce8b4055ceb17f5357ff0e0184ea7b46a5cccb9f46eea3fd3bda7d85236a07a73019728531dbab8fe25f324436b9c3067234ba05fa4cb227e9aa14e436450cf457fa686a82dcd77a0ac6ee3b6f53c0b8d134fe884d9144f0055e83277e5af23471d2bcfd1ff2b64190db0657c6c50c728b59419acbe6d1c669de90ac84ff84ac4135a65e94e86333c15ea43838c666191e08dd2a6c004d8e82665de1914fbfffc49dc55c1ee2a59f89a920e62d03edec78c5ad751dffefefc964e25115911ac4bd1ca93eeefa33da30ed4c7ba7da465bb347bb06a06aa8dfeddb61bae053322e06267510383f903954b4dd522d7c49b58b57fba3b410754edb93f2fd3d50d22dbfba0252ff03a2eb95a66ce5a9edbae958852af0e014f378880847844bc75d57f9d1cb624126e90c0cdd8f1022ff447733bb8ecc1cd35eb13f6d41bb89106cba5eddee177f234f717c36dea9edcdeeac034e991cb64e25235bf6c2b70ec0a463134688150a9fe9412395c37608a43558c96b1a86a4c8745ce7383b95afa00457599dd3092a13c49111501e9d24c9d4754a47f36245e3478afab05096d1ac3812f7f8b0161c018d78429a2468be49c2a6321c694d4a369c154ba8e7838925f8e7aa61325435646d8df4ac3cbec7802a83b7a9085699794bdc43b524c9365e6e2fd3ecade9f33db5d4fd11fe196dabb18bb10097c86653ae8beee5a306bb6f68169b8720649cd12bf190833d596f4828c9de3ec40d1287679c4c9b0be933ee267272b9aa8fcec6a9840b7072fd6c4926b5ba381ab53562a27d2223d63a14ee12076bdd70ae5d21620ac7eec86163aa8011781fcb6913db666522f72e248028aae33d79da2d6417d7dce294769fcb8fb597e005cbd3756c3cee68c761bccd2e56402498e9185a10be580c621aa82a72c2b79c17589f2ebda0c9a8b841145f74eb1998b16706c86abd7e44f1b2272ac0ede829921f91f87775e970f2df654c22d3f0773037a166e86d6cfe85d5b33aba771f274aa079c2647d9c256e74a53b1fdda30d85c169deb45616e4929d51b7725e66331cdf05c4f6ca757e2d3ca4369efb9b38d9fffefc3c3f8dbf8a2a9e8106902c12957336173097367a4b9187df3df50398c2ef414ca13dd5b8bb998d2d21c8c94d44c523978ac7de8d63039b2e28f7fc621360655522b4d98fe4bbe4956c1da3ae03ff16179310dd37e1254182ab8c183311aa13abb2e30c4b4aa33316f00e8414fc760b3bd8c9433bc8585615343eebf966325378a3c73187d70563f5914d476fb3eb3971c7cf26d9551c5ad40b44b6f78b9538778c92de3e513361ff9584eb2345d9fd60448994f07f5f0b454ac7feef9ba5a6ebf6540133c7a7a88bef5433abb7449f42a21f7701694eea0f61bdec567ee3e19615b78c38ab8ce1f7af0223dad7fed526f7dddc6fba11f61090eaddf91d90ee772c2bbcb9dae54361389978eecc113e106e57e0cc9638429bad9fc570d50cb481bc478b6b073fcb76651ee661904635ea4b5f645ee5aea1fd1331c7e7aa1657067da4201a933fae899863affba0f581e0ed17a7095ed40191707ad2f89d3b677f33557b5d0fbb358d38adf0a7cac5589415a2c6103cf08724e15f20c0810cb3e0821d359f69cf1d2cf581797f291b7e34d427cf3bce9194533af8fa401448e87ec391782662a921dd316d4f06a7c29d19f82ca3621b0867c6b430158859b3a9070f955fa41c71c8cca3f63f2f6d9bbb38075ac63eabd3cde4323e5dc3cf7a572fcffadabb65f790ac3650d67d307457f38ec662176ffdb41ccab76b039ef1f082cd562d594cb0fce7edd73cceef9bd8ffa35aa1f91ee3052c01d35bcc14b41e06b3af5053bfe58525a70d5c369ec3c2c3627cdc342f02b5b3bef42f9a0f2eef063f74b0df9bc5c845b4ecb0f37eb93888dbda61a7afd298909e6c3af8e8ee01d9abdc33382474ea1f38eb7b9a8d312bb3067cbac7abb72be64af5fc70b0a244dd922eb9cfbcb4d4b438f8cf58b3b463f6e95af0b669c3790b433f4406ff0aafccca93761f23941ff5306e860bc536a7e9f875aae979869b8de55ab696f6a51f05daaeecd18c3c22b9e398412025864828389e2f4ff0e195d62acd32f5090ee1a8e9f0243565a758ad3f46aa0b3cbeef25584a1ae0017222f393d4e4f53b300000000000000000000000000000000000000000000000000090f13161e242832;
                             
              
        #140;

        $finish;
    end
    
    always begin 
    #0.001 clk = ~clk;
    end

    // Dump waveforms for debugging
    initial begin
        $dumpfile("verifyTop_tb.vcd");
        $dumpvars(0, verifyTop_tb);
    end
endmodule