module Chi(
    input  logic [63:0] A [0:4][0:4],  // 64-bit elements in a 5x5 matrix
    output logic [63:0] Ab[0:4][0:4]   // 64-bit output elements in a 5x5 matrix
);

    // Static, explicit computation for each matrix element

    // Row 0
    always_comb begin
    Ab[0][0] = A[0][0]^(~A[1][0]&A[2][0]);
    Ab[0][1] = A[0][1] ^ (~A[1][1] & A[2][1]);
    Ab[0][2] = A[0][2] ^ (~A[1][2] & A[2][2]);
    Ab[0][3] = A[0][3] ^ (~A[1][3] & A[2][3]);
    Ab[0][4] = A[0][4] ^ (~A[1][4] & A[2][4]);

    // Row 1
    Ab[1][0] = A[1][0] ^ (~A[2][0] & A[3][0]);
    Ab[1][1] = A[1][1] ^ (~A[2][1] & A[3][1]);
    Ab[1][2] = A[1][2] ^ (~A[2][2] & A[3][2]);
    Ab[1][3] = A[1][3] ^ (~A[2][3] & A[3][3]);
    Ab[1][4] = A[1][4] ^ (~A[2][4] & A[3][4]);

    // Row 2
    Ab[2][0] = A[2][0] ^ (~A[3][0] & A[4][0]);
    Ab[2][1] = A[2][1] ^ (~A[3][1] & A[4][1]);
    Ab[2][2] = A[2][2] ^ (~A[3][2] & A[4][2]);
    Ab[2][3] = A[2][3] ^ (~A[3][3] & A[4][3]);
    Ab[2][4] = A[2][4] ^ (~A[3][4] & A[4][4]);

    // Row 3
    Ab[3][0] = A[3][0] ^ (~A[4][0] & A[0][0]);
    Ab[3][1] = A[3][1] ^ (~A[4][1] & A[0][1]);
    Ab[3][2] = A[3][2] ^ (~A[4][2] & A[0][2]);
    Ab[3][3] = A[3][3] ^ (~A[4][3] & A[0][3]);
    Ab[3][4] = A[3][4] ^ (~A[4][4] & A[0][4]);

    // Row 4
    Ab[4][0] = A[4][0] ^ (~A[0][0] & A[1][0]);
    Ab[4][1] = A[4][1] ^ (~A[0][1] & A[1][1]);
    Ab[4][2] = A[4][2] ^ (~A[0][2] & A[1][2]);
    Ab[4][3] = A[4][3] ^ (~A[0][3] & A[1][3]);
    Ab[4][4] = A[4][4] ^ (~A[0][4] & A[1][4]);
    end


   
endmodule
